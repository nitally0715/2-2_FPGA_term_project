//==============================================================
// Money_Manager.v (FINAL Version - port name unified)
// - FSM_Controller / Hit_Check / Top_Roulette�� ���� ����
//==============================================================

module Money_Manager(
    input  wire        clk,
    input  wire        rst,

    // FSM �� Money_Manager
    input  wire        update_req,     // �ܾ� ���� ��û (1Ŭ��)
    input  wire        win_flag,       // Hit_Check ��� (��/��)  <-- �̸� ����!
    input  wire [15:0] bet_amount,     // ���� �ݾ�
    input  wire [2:0]  bet_count,      // ���� ����(1~4)
    input  wire [2:0]  hit_count,      // ���� ����

    // Money_Manager �� FSM / Display / Top
    output reg [15:0] current_money,   // ���� �ܾ� (0~10000)
    output reg        money_zero,      // �ܾ� == 0
    output reg        money_10000,     // �ܾ� >= 10000 (���� Ŭ����)
    output reg        win_flag_out     // FSM ���޿� �н�����
);

    //==========================================================
    // �ʱ� �ں�
    //==========================================================
    localparam INITIAL_MONEY = 16'd100;
    localparam MAX_MONEY     = 16'd10000;

    //==========================================================
    // ��� ��� ��� : bet_count�� ���� payout ��� ����
    //==========================================================
    reg [3:0] payout_multi;

    always @(*) begin
        case (bet_count)
            3'd1: payout_multi = 4'd8;
            3'd2: payout_multi = 4'd4;
            3'd3: payout_multi = 4'd2;
            3'd4: payout_multi = 4'd1;
            default: payout_multi = 4'd0;
        endcase
    end

    //==========================================================
    // update_req rising-edge detect
    //==========================================================
    reg update_req_prev;
    wire update_pulse = (update_req == 1'b1 && update_req_prev == 1'b0);

    always @(posedge clk or posedge rst) begin
        if (rst)
            update_req_prev <= 1'b0;
        else
            update_req_prev <= update_req;
    end

    //==========================================================
    // ���� �ӽ� ��������
    //==========================================================
    reg [31:0] payout;
    reg [31:0] temp_money;

    //==========================================================
    // Money Update Logic
    //==========================================================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            current_money <= INITIAL_MONEY;
            money_zero    <= 1'b0;
            money_10000   <= 1'b0;
            win_flag_out  <= 1'b0;
        end else begin
            // Hit_Check �� FSM �� Money_Manager �н� ����
            win_flag_out <= win_flag;

            //------------------------------------------------------
            // update_req 1Ŭ�� �� �ܾ� ����
            //------------------------------------------------------
            if (update_pulse) begin

                // �й�
                if (!win_flag) begin
                    if (current_money > bet_amount)
                        current_money <= current_money - bet_amount;
                    else
                        current_money <= 16'd0;
                end

                // �¸�
                else begin
                    payout = bet_amount * payout_multi;

                    temp_money = current_money;

                    // ���ñ� ����
                    if (temp_money > bet_amount)
                        temp_money = temp_money - bet_amount;
                    else
                        temp_money = 0;

                    // ���� ����
                    temp_money = temp_money + payout;

                    // ���� ����
                    if (temp_money >= MAX_MONEY)
                        current_money <= MAX_MONEY;
                    else
                        current_money <= temp_money[15:0];
                end
            end

            //------------------------------------------------------
            // �ܾ� ���� �÷��� ������Ʈ
            //------------------------------------------------------
            money_zero  <= (current_money == 16'd0);
            money_10000 <= (current_money >= MAX_MONEY);
        end
    end

endmodule
