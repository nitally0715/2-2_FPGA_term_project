//==============================================================
// Roulette_LED.v
// - 8���� LED�� �̿��� �귿 ȸ��/����/���� ǥ��
// - FSM_Controller �� start_spin(1Ŭ��) �Է��� �޾� ����
// - ��� ��ġ result_pos(0~7) ���
// - LFSR�� �̿��ؼ� ������ �ο�
//==============================================================

module Roulette_LED(
    input  wire clk,
    input  wire rst,
    input  wire start_spin,       // FSM���� 1Ŭ�� �޽�

    output reg  [7:0] led_out,    // ���� LED ��� (one-hot)
    output reg  [2:0] result_pos, // ���� ���� ��ġ (0~7)
    output reg        spin_done,  // ȸ�� ���� ��ȣ (1Ŭ�� �޽�)
    output reg        spin_active // ȸ�� ���� �� 1 (RUN, SLOW ����)
);

    //==========================================================
    // 0. ȸ�� FSM ���� ����
    //==========================================================
    localparam  S_IDLE = 2'd0,
                S_RUN  = 2'd1,
                S_SLOW = 2'd2,
                S_STOP = 2'd3;

    reg [1:0] state, state_next;

    //==========================================================
    // 1. ���� pos (0~7)
    //==========================================================
    reg [2:0] pos;  // ���� LED �ε���

    // LED one-hot ���� (active-high)
    wire [7:0] led_pattern = (8'b0000_0001 << pos);

    //==========================================================
    // 2. �ӵ� ����� ���ֱ�
    //==========================================================
    reg [31:0] speed_cnt;
    reg [31:0] interval;       // ���� ������ (�������� ����)

    // ��� ȸ�� �⺻�ӵ� & ���� ������
    localparam BASE_SPEED   = 32'd2_000_000;   // 50MHz ���� �� 40ms
    localparam SLOW_STEP    = 32'd200_000;     // ���� �ܰ� ������
    localparam MAX_INTERVAL = 32'd12_000_000;  // ���� �Ѱ�

    //==========================================================
    // 3. LFSR(���� ����)
    //==========================================================
    reg [7:0] lfsr;

    always @(posedge clk or posedge rst) begin
        if (rst)
            lfsr <= 8'hA5; // �ʱ� seed
        else begin
            // x^8 + x^6 + x^5 + x^4 + 1 ���׽�
            lfsr <= {lfsr[6:0], lfsr[7] ^ lfsr[5] ^ lfsr[4] ^ lfsr[3]};
        end
    end

    //==========================================================
    // 4. ���� ��������
    //==========================================================
    always @(posedge clk or posedge rst) begin
        if (rst)
            state <= S_IDLE;
        else
            state <= state_next;
    end

    //==========================================================
    // 5. ���� ���� ���� (���� ��)
//==========================================================
    always @(*) begin
        state_next = state;
        case (state)
            //--------------------------------------------------
            // IDLE
            //--------------------------------------------------
            S_IDLE: begin
                if (start_spin)
                    state_next = S_RUN;
            end

            //--------------------------------------------------
            // ��� ȸ��
            //--------------------------------------------------
            S_RUN: begin
                // interval�� ���� ���� �̻� Ŀ���� ���� �ܰ��
                if (interval >= (BASE_SPEED + SLOW_STEP * 4))
                    state_next = S_SLOW;
            end

            //--------------------------------------------------
            // ���� ��
            //--------------------------------------------------
            S_SLOW: begin
                if (interval >= MAX_INTERVAL)
                    state_next = S_STOP;
            end

            //--------------------------------------------------
            // ����
            //--------------------------------------------------
            S_STOP: begin
                // spin_done 1Ŭ�� �� IDLE ����
                state_next = S_IDLE;
            end

            default: begin
                state_next = S_IDLE;
            end
        endcase
    end

    //==========================================================
    // 6. �ӵ� ���� & pos ������Ʈ & ���
    //==========================================================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            pos        <= 3'd0;
            speed_cnt  <= 32'd0;
            interval   <= BASE_SPEED;
            led_out    <= 8'd0;
            result_pos <= 3'd0;
            spin_done  <= 1'b0;
            spin_active<= 1'b0;
        end else begin
            // �⺻��
            led_out     <= led_pattern; // ���� pos ���� one-hot
            spin_done   <= 1'b0;        // �޽� ��ȣ
            spin_active <= 1'b0;        // �⺻�� 0

            case (state)
                //--------------------------------------------------
                // IDLE
                //--------------------------------------------------
                S_IDLE: begin
                    // ���� ���� �� �ӵ� ���� �� �ʱ�ȭ
                    interval  <= BASE_SPEED;
                    speed_cnt <= 32'd0;
                    // LED�� ���� ���� ������ �Ʒ� �ּ��� ����
                    // led_out   <= 8'd0;

                    if (start_spin) begin
                        // ���� ���� ��ġ
                        pos <= lfsr[2:0];
                    end
                end

                //--------------------------------------------------
                // RUN (������ ȸ��)
                //--------------------------------------------------
                S_RUN: begin
                    spin_active <= 1'b1;

                    if (speed_cnt >= interval) begin
                        speed_cnt <= 32'd0;
                        pos       <= pos + 3'd1;  // 0~7 ��ȯ

                        // ������ ���� ����
                        if (interval < (BASE_SPEED + SLOW_STEP * 4))
                            interval <= interval + SLOW_STEP;
                    end else begin
                        speed_cnt <= speed_cnt + 32'd1;
                    end
                end

                //--------------------------------------------------
                // SLOW_DOWN (������ ȸ��)
                //--------------------------------------------------
                S_SLOW: begin
                    spin_active <= 1'b1;

                    if (speed_cnt >= interval) begin
                        speed_cnt <= 32'd0;
                        pos       <= pos + 3'd1;

                        // �� �ް��� ����
                        if (interval < MAX_INTERVAL)
                            interval <= interval + (SLOW_STEP << 1);
                    end else begin
                        speed_cnt <= speed_cnt + 32'd1;
                    end
                end

                //--------------------------------------------------
                // STOP_RESULT
                //--------------------------------------------------
                S_STOP: begin
                    // ���� ��ġ Ȯ��
                    result_pos <= pos;
                    spin_done  <= 1'b1;   // FSM�� ȸ�� ���� �˸� (1Ŭ��)
                    // led_out �� led_pattern���� ���� pos ����
                end

                default: begin
                    // ������
                end
            endcase
        end
    end

endmodule
