//=======================================================================
// Roulette_LED.v  (�ε巯�� ���� + ��Ȯ ���� �ϼ���)
//=======================================================================
module Roulette_LED(
    input  wire clk,          // 50 MHz
    input  wire rst,
    input  wire start,        // FSM�� 1Ŭ�� �޽� ����
    output reg  [7:0] led,    // LED 8�� (active high)
    output reg  [2:0] pos,    // 0~7, ��÷ ��ġ
    output reg  spin_done     // 1Ŭ�� �޽�
);

    //-------------------------------------------------------------
    // ���� ���� ����
    //-------------------------------------------------------------
    reg spinning;             // ȸ�� �� ����
    reg [31:0] delay_cnt;     // ȸ�� �ӵ� ī����
    reg [31:0] delay_max;     // ī��Ʈ ��ǥ�� (���� ����)
    reg [31:0] decel_step;    // ���� ����

    localparam DELAY_FAST  = 32'd200000;   // �ʱ� �ӵ� (����)
    localparam DELAY_SLOW  = 32'd5000000;  // ���� ���� (���߱� ����)
    localparam DECEL_INIT  = 32'd20000;    // ���� �⺻ ������


    //-------------------------------------------------------------
    // ���� �귿 ȸ�� ����
    //-------------------------------------------------------------
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            spinning   <= 0;
            pos        <= 0;
            delay_cnt  <= 0;
            delay_max  <= DELAY_FAST;
            decel_step <= DECEL_INIT;
            spin_done  <= 0;
        end 
        else begin
            spin_done <= 0;

            // ----------------------------------------------------
            // START ��ȣ �� ȸ�� ����
            // ----------------------------------------------------
            if (start && !spinning) begin
                spinning   <= 1;
                delay_max  <= DELAY_FAST;
                decel_step <= DECEL_INIT;
                delay_cnt  <= 0;
            end

            // ----------------------------------------------------
            // ȸ�� ��
            // ----------------------------------------------------
            if (spinning) begin

                // delay_cnt�� delay_max�� �ʰ��ϸ� pos ����
                if (delay_cnt >= delay_max) begin
                    delay_cnt <= 0;

                    // LED ��ġ �� ĭ �̵�
                    pos <= (pos == 3'd7) ? 3'd0 : pos + 1'b1;

                    // ����: ���� delay_max�� Ŀ���� ȸ���� ������
                    if (delay_max < DELAY_SLOW)
                        delay_max <= delay_max + decel_step;
                    else begin
                        // ���� �� �� ����
                        spinning  <= 0;
                        spin_done <= 1;
                    end

                end else begin
                    delay_cnt <= delay_cnt + 1;
                end
            end
        end
    end

    //-------------------------------------------------------------
    // LED ���� ���� (pos ��ġ�� ����)
    //-------------------------------------------------------------
    always @(*) begin
        led = 8'b00000000;
        led[pos] = 1'b1;
    end

endmodule
