//===========================================================
// Piezo_Buzzer.v
// - FSM ���¿� ���� �ٸ� ��/��ε� ���
// - START_SPIN: ���� �ݺ���
// - SPIN_WAIT: ���� �ݺ���
// - WIN_DISPLAY: ª�� ��ε�
// - LOSE_DISPLAY: ���� �����
//===========================================================

module Piezo_Buzzer(
    input  wire clk,          // 50MHz ����
    input  wire rst,
    input  wire [3:0] state,
    output reg  piezo
);

    //----------------------------------------------------
    // �����ڵ�(FSM�� �ݵ�� ��ġ)
    //----------------------------------------------------
    localparam S_START_SPIN   = 4'd4;
    localparam S_SPIN_WAIT    = 4'd5;
    localparam S_WIN_DISPLAY  = 4'd7;
    localparam S_LOSE_DISPLAY = 4'd8;

    //----------------------------------------------------
    // Piezo�� �ܼ� square wave �� divider�� �� ����
    //----------------------------------------------------
    reg [31:0] cnt;
    reg [31:0] tone_div;   // ���ļ� ����
    reg        enable;     // Piezo on/off

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            cnt   <= 0;
            piezo <= 0;
            enable <= 0;
            tone_div <= 32'd0;
        end else begin

            //------------------------------------------------
            // ���º� �� ����
            //------------------------------------------------
            case (state)

                // --------------------------------------------
                // 1) ȸ�� ���� �� ���� 4kHz ������
                // --------------------------------------------
                S_START_SPIN: begin
                    enable   <= 1;
                    tone_div <= 32'd6250;  // 50MHz / 6250 = 8kHz �� /2 �� �� 4kHz
                end

                // --------------------------------------------
                // 2) SPIN_WAIT �� ���� ���� 2.5~3kHz (�߰� �ӵ�)
                // --------------------------------------------
                S_SPIN_WAIT: begin
                    enable   <= 1;
                    tone_div <= 32'd10000; // ~2.5kHz
                end

                // --------------------------------------------
                // 3) �¸� ��ε� (C �� E �� G �� C)
                // --------------------------------------------
                S_WIN_DISPLAY: begin
                    enable <= 1;

                    // ��ε� ����� ī����
                    case (cnt[18:16])   // �� 150ms ����
                        3'd0: tone_div <= 32'd38220; // C (261 Hz)
                        3'd1: tone_div <= 32'd30337; // E (329 Hz)
                        3'd2: tone_div <= 32'd25510; // G (392 Hz)
                        3'd3: tone_div <= 32'd38220; // C (261 Hz)
                        default: tone_div <= 32'd38220;
                    endcase
                end

                // --------------------------------------------
                // 4) �й� �� ���� ����� 300Hz
                // --------------------------------------------
                S_LOSE_DISPLAY: begin
                    enable   <= 1;
                    tone_div <= 32'd41666; // 300Hz
                end

                // --------------------------------------------
                // 5) �� �� = ����
                // --------------------------------------------
                default: begin
                    enable   <= 0;
                    tone_div <= 32'd0;
                end
            endcase


            //------------------------------------------------
            // Tone ���� (Square Wave)
            //------------------------------------------------
            if (enable && tone_div != 0) begin
                cnt <= cnt + 1;
                if (cnt >= tone_div) begin
                    cnt   <= 0;
                    piezo <= ~piezo; // square wave
                end
            end else begin
                cnt   <= 0;
                piezo <= 0;
            end
        end
    end

endmodule
