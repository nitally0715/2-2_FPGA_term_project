//====================================================
// Money_Manager.v
// - ���� �ݾ� / ��� / ���п� ���� �ܾ� ����
// - UPDATE_MONEY ���� �� 1Ŭ�������� ����
//====================================================

module Money_Manager(
    input  wire        clk,
    input  wire        rst,

    input  wire [3:0]  state,        // FSM ����
    input  wire [15:0] bet_amount,   // �Էµ� ���� �ݾ�
    input  wire [2:0]  bet_count,    // �Էµ� ���� ���� (1~4)
    input  wire        win_flag,     // ���� STOP_RESULT���� ������

    output reg [15:0]  current_money // ���� �ܾ�
);

    // FSM ���� ���� (FSM_Controller�� �ݵ�� ��ġ�� ��)
    localparam S_UPDATE_MONEY = 4'd9;
    localparam START_MONEY    = 16'd100;

    // UPDATE_MONEY�� 1ȸ�� �����ϱ� ���� ���� ���� ����
    reg [3:0] prev_state;

    // ��� ��� ���̺� �Լ�
    function [15:0] payout_multiplier(input [2:0] count);
        begin
            case (count)
                1: payout_multiplier = 16'd8;  
                2: payout_multiplier = 16'd4;
                3: payout_multiplier = 16'd3;
                4: payout_multiplier = 16'd2;
                default: payout_multiplier = 16'd1;
            endcase
        end
    endfunction

    //====================================================
    // ���� ����
    //====================================================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            current_money <= START_MONEY;
            prev_state    <= 4'd0;
        end else begin
            prev_state <= state;

            //------------------------------------------------------
            // UPDATE_MONEY ���¿��� "state�� ó�� ������ ��" �� 1ȸ ó��
            //------------------------------------------------------
            if (state == S_UPDATE_MONEY && prev_state != S_UPDATE_MONEY) begin
                
                // ������ġ: ���� �ݾ��� �����ݾ׺��� ���ٸ� ����
                if (bet_amount > current_money) begin
                    // ��� FSM���� �̹� �ݾ� ���������� �����ϰ� ����
                    current_money <= current_money;
                end 
                else if (win_flag) begin
                    // WIN: �߰� ���� = bet_amount * (��� - 1)
                    current_money <= current_money 
                                   + bet_amount * payout_multiplier(bet_count)
                                   - bet_amount;
                end 
                else begin
                    // LOSE: bet_amount��ŭ ����
                    if (current_money > bet_amount)
                        current_money <= current_money - bet_amount;
                    else
                        current_money <= 16'd0;  // 0 �Ʒ��δ� �ȳ�����
                end

            end
        end
    end

endmodule
