//======================================================================
// Piezo_Buzzer.v (50MHz)
// - FSM state / spin_active �� ���� ȿ���� & ��ε� ���
//   * START_SPIN, SLOW_DOWN : ȸ�� ȿ����
//   * WIN_DISPLAY          : ª�� �¸� ��ε� (���ֵ��ٵ�)
//   * LOSE_DISPLAY         : ���� �й���
//   * GAME_CLEAR           : ���� ������ Ŭ���� ���� 4��
//   * ������ ����          : ����
//======================================================================

module Piezo_Buzzer(
    input  wire       clk,         // 50MHz
    input  wire       rst,
    input  wire [3:0] state,
    input  wire       spin_active, // �귿 ȸ�� ���̸� 1
    input  wire       win_flag,    // (������ �� �ᵵ ��, ��Ʈ�� ����)

    output reg        piezo_out
);

    // FSM �����ڵ� (FSM_Controller�� ����� ��)
    localparam S_IDLE         = 4'd0;
    localparam S_BET_MONEY    = 4'd1;
    localparam S_BET_SELECT   = 4'd2;
    localparam S_NUMBER_INPUT = 4'd3;
    localparam S_START_SPIN   = 4'd4;
    localparam S_SLOW_DOWN    = 4'd5;
    localparam S_STOP_RESULT  = 4'd6;
    localparam S_WIN_DISPLAY  = 4'd7;
    localparam S_LOSE_DISPLAY = 4'd8;
    localparam S_UPDATE_MONEY = 4'd9;
    localparam S_CHECK_MONEY  = 4'd10;
    localparam S_NEXT_STAGE   = 4'd11;
    localparam S_GAME_OVER    = 4'd12;
    localparam S_GAME_CLEAR   = 4'd13;

    //==========================================================
    // 1) ��ε�� free-running ī����
    //    -> ���� ��Ʈ�� �߶� "�� ��° ������"�� ���
    //==========================================================
    reg [23:0] mel_cnt;
    always @(posedge clk or posedge rst) begin
        if (rst)
            mel_cnt <= 24'd0;
        else
            mel_cnt <= mel_cnt + 24'd1;
    end

    //==========================================================
    // 2) �� ���ֱ� : 50MHz -> ���ϴ� ���ļ��� �簢��
    //
    //    tone_divider = 0 : ����
    //    tone_divider > 0 : clk�� ������ tone_clk ����
    //
    //    �뷫���� ���ļ� (50MHz ����)
    //      25000 -> �� 1kHz
    //      20000 -> �� 1.25kHz
    //      15000 -> �� 1.6kHz
    //      10000 -> �� 2.5kHz
    //      50000 -> �� 500Hz
    //==========================================================
    reg [31:0] tone_divider;
    reg [31:0] tone_cnt;
    reg        tone_clk;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            tone_cnt  <= 32'd0;
            tone_clk  <= 1'b0;
        end else begin
            if (tone_divider == 32'd0) begin
                // ������ ���� ī���� ���� + ��� 0
                tone_cnt <= 32'd0;
                tone_clk <= 1'b0;
            end else begin
                if (tone_cnt >= tone_divider) begin
                    tone_cnt <= 32'd0;
                    tone_clk <= ~tone_clk;
                end else begin
                    tone_cnt <= tone_cnt + 32'd1;
                end
            end
        end
    end

    //==========================================================
    // 3) ���º� tone_divider ����
    //==========================================================
    always @(*) begin
        // �⺻�� : ����
        tone_divider = 32'd0;

        case (state)

            //--------------------------------------------------
            // ȸ�� ȿ���� : START_SPIN / SLOW_DOWN + spin_active
            //--------------------------------------------------
            S_START_SPIN,
            S_SLOW_DOWN: begin
                if (spin_active) begin
                    // mel_cnt �Ϻ� ��Ʈ�� �ణ�� "��������" ����
                    case (mel_cnt[18:17])
                        2'd0: tone_divider = 32'd22000; // �� 1.1kHz
                        2'd1: tone_divider = 32'd18000; // �� 1.4kHz
                        2'd2: tone_divider = 32'd15000; // �� 1.6kHz
                        default: tone_divider = 32'd18000;
                    endcase
                end else begin
                    tone_divider = 32'd0; // ȸ�� �� �ϸ� ����
                end
            end

            //--------------------------------------------------
            // WIN_DISPLAY : ª�� �¸� ��ε� (���ֵ��ٵ�)
            //--------------------------------------------------
            S_WIN_DISPLAY: begin
                case (mel_cnt[20:19])   // 4�ܰ� �ݺ� (note�� �� ���� ms)
                    2'd0: tone_divider = 32'd20000; // �߰���
                    2'd1: tone_divider = 32'd15000; // �� �� ���� ��
                    2'd2: tone_divider = 32'd20000; // �߰���
                    2'd3: tone_divider = 32'd25000; // �ణ ���� ��
                    default: tone_divider = 32'd0;
                endcase
            end

            //--------------------------------------------------
            // LOSE_DISPLAY : ���� �й��� (��-)
            //--------------------------------------------------
            S_LOSE_DISPLAY: begin
                tone_divider = 32'd50000; // �� 500Hz, ���� ��
            end

            //--------------------------------------------------
            // GAME_CLEAR : ���� 4�� (A-B-A-G ����)
            //--------------------------------------------------
            S_GAME_CLEAR: begin
                case (mel_cnt[21:19])   // 8�ܰ� �� ���� 4�ܰ� ���
                    3'd0: tone_divider = 32'd17000; // A
                    3'd1: tone_divider = 32'd15000; // B (���� ����)
                    3'd2: tone_divider = 32'd17000; // A
                    3'd3: tone_divider = 32'd22000; // G (���� ����)
                    default: tone_divider = 32'd0;
                endcase
            end

            //--------------------------------------------------
            // GAME_OVER : ���� ���� �����
            //--------------------------------------------------
            S_GAME_OVER: begin
                tone_divider = 32'd80000; // �� ���� ��
            end

            //--------------------------------------------------
            // ������ ���� : ����
            //--------------------------------------------------
            default: begin
                tone_divider = 32'd0;
            end
        endcase
    end

    //==========================================================
    // 4) ���� piezo ���
    //==========================================================
    always @(posedge clk or posedge rst) begin
        if (rst)
            piezo_out <= 1'b0;
        else begin
            if (tone_divider == 32'd0)
                piezo_out <= 1'b0;   // ����
            else
                piezo_out <= tone_clk; // �簢�� ���
        end
    end

endmodule
