//====================================================
// FSM_Controller.v
//  - Ű�е� �Է����� ���� �ݾ�/����/��ȣ ����
//  - �귿 ���� ��ȣ(start_spin) �߻�
//  - spin_done ���� ��÷ ���� ����
//  - Money_Manager�� �� win_flag / lose_flag / bet_amount / bet_count ���
//====================================================
module FSM_Controller(
    input  wire        clk,
    input  wire        rst,

    input  wire        key_valid,
    input  wire [3:0]  key_value,      // 0~9, 10='*', 11='#'

    input  wire        spin_done,
    input  wire [2:0]  roulette_pos,   // 0~7 (=> 1~8)
    input  wire [15:0] current_money,  // ���� �ܾ� (Money_Manager ���)

    output reg         start_spin,     // Roulette_LED ���� Ʈ���� (1Ŭ��)
    output reg         win_flag,
    output reg         lose_flag,

    output reg [15:0]  bet_amount,
    output reg [2:0]   bet_count,

    output reg [3:0]   state
);

    //------------------------------------------------
    // ���� ����
    //------------------------------------------------
    localparam S_IDLE         = 4'd0,
               S_BET_AMOUNT   = 4'd1,
               S_BET_COUNT    = 4'd2,
               S_NUM_INPUT    = 4'd3,
               S_START_SPIN   = 4'd4,
               S_SPIN_WAIT    = 4'd5,
               S_STOP_RESULT  = 4'd6,
               S_WIN_DISPLAY  = 4'd7,
               S_LOSE_DISPLAY = 4'd8,
               S_UPDATE_MONEY = 4'd9,
               S_CHECK_OVER   = 4'd10,
               S_GAME_OVER    = 4'd11;

    //------------------------------------------------
    // ���� �����: ���� ��ȣ �ִ� 4��
    //------------------------------------------------
    reg [3:0] bet_nums [0:3];    // 1~8 ����
    reg [2:0] num_idx;           // �� �� �Է��ߴ���

    // ��� ��ȣ (1~8)
    wire [3:0] result_num = roulette_pos + 1;

    // ���÷��̿� ���� �ð� ī���� (WIN/LOSE ���� ����)
    reg [15:0] disp_cnt;

    // for-loop�� ������ ��� ��ܿ� ����
    integer i;


    //------------------------------------------------
    // ���� FSM
    //------------------------------------------------
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state      <= S_IDLE;
            bet_amount <= 16'd0;
            bet_count  <= 3'd0;
            num_idx    <= 3'd0;
            start_spin <= 1'b0;
            win_flag   <= 1'b0;
            lose_flag  <= 1'b0;
            disp_cnt   <= 16'd0;
        end else begin
            // �⺻��
            start_spin <= 1'b0;

            case (state)

                //------------------------------------------------
                // 0. ��� ����
                //------------------------------------------------
                S_IDLE: begin
                    bet_amount <= 16'd0;
                    bet_count  <= 3'd0;
                    num_idx    <= 3'd0;
                    win_flag   <= 1'b0;
                    lose_flag  <= 1'b0;

                    // '*' �� ���� ���� (�ܾ� > 0 �� ����)
                    if (key_valid && key_value == 4'd10 && current_money > 0)
                        state <= S_BET_AMOUNT;
                end

                //------------------------------------------------
                // 1. ���� �ݾ� �Է� (���� ������ '*' Ȯ��, '#' �ʱ�ȭ)
                //------------------------------------------------
                S_BET_AMOUNT: begin
                    if (key_valid) begin
                        if (key_value <= 4'd9) begin
                            // 10���� �ڸ��� �߰�
                            bet_amount <= bet_amount * 10 + key_value;
                        end else if (key_value == 4'd11) begin
                            // '#': �ٽ� �Է�
                            bet_amount <= 16'd0;
                        end else if (key_value == 4'd10) begin
                            // '*': Ȯ�� (0���� ũ��, �ܾ� ������ ����)
                            if (bet_amount > 0 && bet_amount <= current_money)
                                state <= S_BET_COUNT;
                        end
                    end
                end

                //------------------------------------------------
                // 2. ���� ����(1~4) �Է�
                //------------------------------------------------
                S_BET_COUNT: begin
                    if (key_valid) begin
                        if (key_value >= 4'd1 && key_value <= 4'd4) begin
                            bet_count <= key_value[2:0];
                            num_idx   <= 3'd0;
                            state     <= S_NUM_INPUT;
                        end else if (key_value == 4'd11) begin
                            // '#': �ݾ� �ܰ�� ���ư���
                            state <= S_BET_AMOUNT;
                        end
                    end
                end

                //------------------------------------------------
                // 3. ��ȣ �Է� (1~8), bet_count ������ŭ
                //------------------------------------------------
                S_NUM_INPUT: begin
                    if (key_valid) begin
                        if (key_value >= 4'd1 && key_value <= 4'd8) begin
                            // ��ȣ ����
                            bet_nums[num_idx] <= key_value;
                            num_idx <= num_idx + 1'b1;

                            // ������ �������� �Է� �Ϸ������� SPIN����
                            if (num_idx == bet_count - 1)
                                state <= S_START_SPIN;
                        end else if (key_value == 4'd11) begin
                            // '#': ��ȣ ���� �ٽ�
                            num_idx <= 3'd0;
                        end
                    end
                end

                //------------------------------------------------
                // 4. �귿 ȸ�� ���� (start_spin 1Ŭ�� �޽�)
                //------------------------------------------------
                S_START_SPIN: begin
                    start_spin <= 1'b1;
                    state      <= S_SPIN_WAIT;
                end

                //------------------------------------------------
                // 5. spin_done ��ȣ ��ٸ���
                //------------------------------------------------
                S_SPIN_WAIT: begin
                    if (spin_done)
                        state <= S_STOP_RESULT;
                end

                //------------------------------------------------
                // 6. ��� ����
                //------------------------------------------------
                S_STOP_RESULT: begin
                    win_flag  <= 1'b0;
                    lose_flag <= 1'b0;

                    // bet_count ������ŭ�� ��
                    for (i = 0; i < 4; i = i + 1) begin
                        if (i < bet_count && bet_nums[i] == result_num)
                            win_flag <= 1'b1;
                    end

                    // lose_flag�� win_flag�� �ݴ�
                    // (���� Ŭ������ �� �� �����ǰ�, ���� win_flag ���� ��� ��)
                    if (!win_flag)
                        lose_flag <= 1'b1;

                    disp_cnt <= 16'd0;
                    if (win_flag)
                        state <= S_WIN_DISPLAY;
                    else
                        state <= S_LOSE_DISPLAY;
                end

                //------------------------------------------------
                // 7. �¸� �޽��� ��� ����
                //------------------------------------------------
                S_WIN_DISPLAY: begin
                    disp_cnt <= disp_cnt + 1'b1;
                    if (disp_cnt == 16'h0FFF)  // ������ ������
                        state <= S_UPDATE_MONEY;
                end

                //------------------------------------------------
                // 8. �й� �޽��� ��� ����
                //------------------------------------------------
                S_LOSE_DISPLAY: begin
                    disp_cnt <= disp_cnt + 1'b1;
                    if (disp_cnt == 16'h0FFF)
                        state <= S_UPDATE_MONEY;
                end

                //------------------------------------------------
                // 9. �ܾ� ������ Money_Manager �ʿ��� ó��
                //------------------------------------------------
                S_UPDATE_MONEY: begin
                    state <= S_CHECK_OVER;
                end

                //------------------------------------------------
                // 10. Game Over ���� Ȯ��
                //------------------------------------------------
                S_CHECK_OVER: begin
                    if (current_money == 16'd0)
                        state <= S_GAME_OVER;
                    else
                        state <= S_IDLE;
                end

                //------------------------------------------------
                // 11. GAME OVER ���� (�ٽ� ������ �������� ó��)
                //------------------------------------------------
                S_GAME_OVER: begin
                    // ���⼭�� �׳� �ӹ���,
                    // �ʿ��ϸ� key �Է����� IDLE�� ���ư��� ���� ����
                    if (key_valid && key_value == 4'd11) // '#'�� ���� ���� ����
                        state <= S_IDLE;
                end

                default: state <= S_IDLE;

            endcase
        end
    end

endmodule
