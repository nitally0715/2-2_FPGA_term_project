//==============================================================
// FSM_Controller.v  (FINAL / Hit_Check + Money_Manager ���� ����)
// - Keypad / Roulette_LED / Hit_Check / Money_Manager / Display ��ü �帧 ����
//==============================================================

module FSM_Controller(
    input  wire        clk,
    input  wire        rst,

    // Keypad �Է�
    input  wire        key_valid,
    input  wire [3:0]  key_value,      // 0~9, 10='*', 11='#'

    // Roulette & Money �÷���
    input  wire        spin_done,      // Roulette_LED ȸ�� �Ϸ�
    input  wire        win_flag,       // Hit_Check���� ���� �¸� ����
    input  wire        money_zero,     // Money_Manager: �ܾ� == 0
    input  wire        money_10000,    // Money_Manager: �ܾ� >= 10000
    input  wire [15:0] current_money,  // Money_Manager: ���� �ܾ� (BET_MONEY ������)

    // FSM ���
    output reg  [3:0]  state,          // ���� ���� �ڵ� (LCD, Piezo ��� ���)
    output reg  [2:0]  bet_count,      // ���� ����(1~4)
    output reg  [15:0] bet_amount,     // ���� �ݾ�
    output reg         clear_input,    // Ű�е� �Է� ���� �ʱ�ȭ (1Ŭ�� �޽�)
    output reg         start_spin,     // �귿 ���� Ʈ���� (1Ŭ�� �޽�)
    output reg         update_money_req, // �ܾ� ���� ��û (1Ŭ��)
    output reg         reset_round,    // �� ��/���� ���¿� (1Ŭ��)

    // Hit_Check �� ���� ���� ��ȣ 4��
    output reg  [3:0]  user_num0,
    output reg  [3:0]  user_num1,
    output reg  [3:0]  user_num2,
    output reg  [3:0]  user_num3
);

    //==========================================================
    // ���� ���� (�ٸ� ���� �����ϰ� ���� ����� ��)
    //==========================================================
    localparam S_IDLE         = 4'd0;
    localparam S_BET_MONEY    = 4'd1;
    localparam S_BET_SELECT   = 4'd2;
    localparam S_NUMBER_INPUT = 4'd3;
    localparam S_START_SPIN   = 4'd4;
    localparam S_SLOW_DOWN    = 4'd5;
    localparam S_STOP_RESULT  = 4'd6;
    localparam S_WIN_DISPLAY  = 4'd7;
    localparam S_LOSE_DISPLAY = 4'd8;
    localparam S_UPDATE_MONEY = 4'd9;
    localparam S_CHECK_MONEY  = 4'd10;
    localparam S_NEXT_STAGE   = 4'd11;
    localparam S_GAME_OVER    = 4'd12;
    localparam S_GAME_CLEAR   = 4'd13;

    reg [3:0] state_next;
    reg [2:0] numbers_entered;   // NUMBER_INPUT���� ���� �Էµ� ����

    //==========================================================
    // ���� �� : ����, �������� ������Ʈ
    //==========================================================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state            <= S_IDLE;
            bet_amount       <= 16'd0;
            bet_count        <= 3'd0;
            numbers_entered  <= 3'd0;

            clear_input      <= 1'b0;
            start_spin       <= 1'b0;
            update_money_req <= 1'b0;
            reset_round      <= 1'b0;

            // ���� ��ȣ �ʱ�ȭ
            user_num0        <= 4'd0;
            user_num1        <= 4'd0;
            user_num2        <= 4'd0;
            user_num3        <= 4'd0;
        end else begin
            state <= state_next;

            // �޽��� ��ȣ �⺻�� 0
            clear_input      <= 1'b0;
            start_spin       <= 1'b0;
            update_money_req <= 1'b0;
            reset_round      <= 1'b0;

            case (state)

                //--------------------------------------------------
                // IDLE : ��� (PRESS * TO START)
                //--------------------------------------------------
                S_IDLE: begin
                    if (key_valid && key_value == 4'd10) begin // '*'
                        reset_round     <= 1'b1;   // Hit_Check, Money_Manager �� ���� ���� ����
                        bet_amount      <= 16'd0;
                        bet_count       <= 3'd0;
                        numbers_entered <= 3'd0;

                        // ���� ��ȣ �ʱ�ȭ
                        user_num0       <= 4'd0;
                        user_num1       <= 4'd0;
                        user_num2       <= 4'd0;
                        user_num3       <= 4'd0;
                    end
                end

                //--------------------------------------------------
                // BET_MONEY : ���� �ݾ� �Է�
                //--------------------------------------------------
                S_BET_MONEY: begin
                    if (key_valid) begin
                        if (key_value <= 4'd9) begin
                            // 10���� ����: ���� *10 + �� �ڸ�
                            bet_amount <= (bet_amount * 10) + key_value;

                        end else if (key_value == 4'd11) begin
                            // '#' : �ݾ� �ʱ�ȭ
                            bet_amount  <= 16'd0;
                            clear_input <= 1'b1;

                        end else if (key_value == 4'd10) begin
                            // '*' : Ȯ�� �õ� �� �߸��� ���̸� ���⼭ �ٷ� �ʱ�ȭ
                            // �߸��� ���: 0�� �̰ų�, ���� �ں����� ū �ݾ�
                            if (bet_amount == 16'd0 || bet_amount > current_money) begin
                                bet_amount  <= 16'd0;
                                clear_input <= 1'b1;
                            end
                        end
                    end
                end

                //--------------------------------------------------
                // BET_SELECT : ���� ���� (1~4)
                //--------------------------------------------------
                S_BET_SELECT: begin
                    if (key_valid) begin
                        if (key_value >= 4'd1 && key_value <= 4'd4) begin
                            bet_count <= key_value[2:0];

                        end else if (key_value == 4'd11) begin
                            // '#' : ���� �ʱ�ȭ
                            bet_count   <= 3'd0;
                            clear_input <= 1'b1;

                        end else if (key_value == 4'd10) begin
                            // '*' : Ȯ�� �õ� �� �߸��Ǹ� ����
                            if (bet_count < 3'd1 || bet_count > 3'd4) begin
                                bet_count   <= 3'd0;
                                clear_input <= 1'b1;
                            end
                        end
                    end
                end

                //--------------------------------------------------
                // NUMBER_INPUT : ��ȣ �Է� (1~8, bet_count��)
                //--------------------------------------------------
                S_NUMBER_INPUT: begin
                    if (key_valid) begin
                        if (key_value >= 4'd1 && key_value <= 4'd8) begin
                            // ��ȿ ��ȣ �Է� + ���� �� ���� �� ���� ��
                            if (numbers_entered < bet_count) begin
                                case (numbers_entered)
                                    3'd0: user_num0 <= key_value;
                                    3'd1: user_num1 <= key_value;
                                    3'd2: user_num2 <= key_value;
                                    3'd3: user_num3 <= key_value;
                                    default: ; // do nothing
                                endcase
                                numbers_entered <= numbers_entered + 3'd1;
                            end

                        end else if (key_value == 4'd11) begin
                            // '#' : ��ü �ʱ�ȭ
                            numbers_entered <= 3'd0;
                            clear_input     <= 1'b1;

                            user_num0       <= 4'd0;
                            user_num1       <= 4'd0;
                            user_num2       <= 4'd0;
                            user_num3       <= 4'd0;

                        end else if (key_value == 4'd10) begin
                            // '*' : Ȯ�� �õ�
                            if (numbers_entered != bet_count || bet_count == 3'd0) begin
                                numbers_entered <= 3'd0;
                                clear_input     <= 1'b1;

                                user_num0       <= 4'd0;
                                user_num1       <= 4'd0;
                                user_num2       <= 4'd0;
                                user_num3       <= 4'd0;
                            end
                        end
                    end
                end

                //--------------------------------------------------
                // START_SPIN : �귿 ���� Ʈ����
                //--------------------------------------------------
                S_START_SPIN: begin
                    start_spin <= 1'b1;   // 1Ŭ�� �޽� �� Roulette_LED ����
                end

                //--------------------------------------------------
                // S_SLOW_DOWN : �귿 ���� / ȸ�� ��
                //--------------------------------------------------
                S_SLOW_DOWN: begin
                    // spin_done�� ��ٸ��� ���� (Roulette_LED���� �ö��)
                end

                //--------------------------------------------------
                // STOP_RESULT : ��� Ȯ��
                //--------------------------------------------------
                S_STOP_RESULT: begin
                    // Hit_Check�� result_pos ������� win_flag�� ������ ���Ҵٰ� ����
                end

                //--------------------------------------------------
                // WIN_DISPLAY : �¸� �� Money_Manager�� ���� ��û
                //--------------------------------------------------
                S_WIN_DISPLAY: begin
                    update_money_req <= 1'b1;   // 1Ŭ�� �޽�
                end

                //--------------------------------------------------
                // LOSE_DISPLAY : �й� �� Money_Manager�� ���� ��û
                //--------------------------------------------------
                S_LOSE_DISPLAY: begin
                    update_money_req <= 1'b1;   // 1Ŭ�� �޽�
                end

                //--------------------------------------------------
                // UPDATE_MONEY : Money_Manager ���� (��� ���̶�� ����)
                //--------------------------------------------------
                S_UPDATE_MONEY: begin
                    // ���� ���� ����
                end

                //--------------------------------------------------
                // CHECK_MONEY : �ܾ� ���� Ȯ��
                //--------------------------------------------------
                S_CHECK_MONEY: begin
                    // money_zero / money_10000 �� Money_Manager���� ����
                end

                //--------------------------------------------------
                // NEXT_STAGE : ���� ���� ����
                //--------------------------------------------------
                S_NEXT_STAGE: begin
                    if (key_valid && key_value == 4'd10) begin // '*'
                        reset_round     <= 1'b1;   // Hit_Check ��ȣ / ���� ī���� ����
                        bet_amount      <= 16'd0;
                        bet_count       <= 3'd0;
                        numbers_entered <= 3'd0;

                        user_num0       <= 4'd0;
                        user_num1       <= 4'd0;
                        user_num2       <= 4'd0;
                        user_num3       <= 4'd0;
                    end
                end

                //--------------------------------------------------
                // GAME_OVER : �ܾ� 0
                //--------------------------------------------------
                S_GAME_OVER: begin
                    if (key_valid && key_value == 4'd10) begin
                        reset_round     <= 1'b1;
                        bet_amount      <= 16'd0;
                        bet_count       <= 3'd0;
                        numbers_entered <= 3'd0;

                        user_num0       <= 4'd0;
                        user_num1       <= 4'd0;
                        user_num2       <= 4'd0;
                        user_num3       <= 4'd0;
                    end
                end

                //--------------------------------------------------
                // GAME_CLEAR : �ܾ� >= 10000 (���� Ŭ����)
                //--------------------------------------------------
                S_GAME_CLEAR: begin
                    if (key_valid && key_value == 4'd10) begin
                        reset_round     <= 1'b1;
                        bet_amount      <= 16'd0;
                        bet_count       <= 3'd0;
                        numbers_entered <= 3'd0;

                        user_num0       <= 4'd0;
                        user_num1       <= 4'd0;
                        user_num2       <= 4'd0;
                        user_num3       <= 4'd0;
                    end
                end

                default: begin
                    // ������: ���� ó�� ����, state_next�� �˾Ƽ� IDLE�� ���� ��
                end
            endcase
        end
    end

    //==========================================================
    // ���� �� : ���� ���� ����
    //==========================================================
    always @(*) begin
        state_next = state;

        case (state)

            //--------------------------------------------------
            S_IDLE: begin
                if (key_valid && key_value == 4'd10)
                    state_next = S_BET_MONEY;
            end

            //--------------------------------------------------
            S_BET_MONEY: begin
                // '*' ���Ȱ�, bet_amount�� 0�� �ƴϰ� current_money �����̸� BET_SELECT��
                if (key_valid && key_value == 4'd10) begin
                    if (bet_amount != 16'd0 && bet_amount <= current_money)
                        state_next = S_BET_SELECT;
                    else
                        state_next = S_BET_MONEY; // �߸��� �Է� �� �ٽ� BET_MONEY
                end
            end

            //--------------------------------------------------
            S_BET_SELECT: begin
                if (key_valid && key_value == 4'd10) begin
                    if (bet_count >= 3'd1 && bet_count <= 3'd4)
                        state_next = S_NUMBER_INPUT;
                    else
                        state_next = S_BET_SELECT;
                end
            end

            //--------------------------------------------------
            S_NUMBER_INPUT: begin
                if (key_valid && key_value == 4'd10) begin
                    if (numbers_entered == bet_count && bet_count != 3'd0)
                        state_next = S_START_SPIN;
                    else
                        state_next = S_NUMBER_INPUT;
                end
            end

            //--------------------------------------------------
            S_START_SPIN: begin
                state_next = S_SLOW_DOWN;
            end

            //--------------------------------------------------
            S_SLOW_DOWN: begin
                if (spin_done)
                    state_next = S_STOP_RESULT;
            end

            //--------------------------------------------------
            S_STOP_RESULT: begin
                // Hit_Check���� ���� win_flag�� ���� ��/�� �б�
                if (win_flag)
                    state_next = S_WIN_DISPLAY;
                else
                    state_next = S_LOSE_DISPLAY;
            end

            //--------------------------------------------------
            S_WIN_DISPLAY: begin
                state_next = S_UPDATE_MONEY;
            end

            //--------------------------------------------------
            S_LOSE_DISPLAY: begin
                state_next = S_UPDATE_MONEY;
            end

            //--------------------------------------------------
            S_UPDATE_MONEY: begin
                state_next = S_CHECK_MONEY;
            end

            //--------------------------------------------------
            S_CHECK_MONEY: begin
                if (money_zero)
                    state_next = S_GAME_OVER;
                else if (money_10000)
                    state_next = S_GAME_CLEAR;
                else
                    state_next = S_NEXT_STAGE;
            end

            //--------------------------------------------------
            S_NEXT_STAGE: begin
                // '*' ������ ���� ���� �� BET_MONEY
                if (key_valid && key_value == 4'd10)
                    state_next = S_BET_MONEY;
            end

            //--------------------------------------------------
            S_GAME_OVER: begin
                // '*' ������ ���� �ʱ�ȭ �� IDLE
                if (key_valid && key_value == 4'd10)
                    state_next = S_IDLE;
            end

            //--------------------------------------------------
            S_GAME_CLEAR: begin
                // '*' ������ ���� �ʱ�ȭ �� IDLE
                if (key_valid && key_value == 4'd10)
                    state_next = S_IDLE;
            end

            default: begin
                state_next = S_IDLE;
            end
        endcase
    end

endmodule
