//====================================================================
// SevenSegment_Display.v
// 5�ڸ� 7-seg ���÷��� ����
// current_money(0~10000) ǥ��, �ʰ� �� 10000���� ����
// active-low ��� (�Ϲ����� FPGA ���� ����)
//
//====================================================================

module SevenSegment_Display(
    input  wire        clk,
    input  wire        rst,
    input  wire [15:0] current_money,   // 0~10000���� ��ȿ

    output reg  [6:0]  seg,             // active-low 7-seg (a~g)
    output reg  [4:0]  an               // active-low �ڸ� ���� 5�ڸ�
);

    //============================================================
    // ���� �� Ŭ����: 0~10000�� ���
    //============================================================
    reg [15:0] money_clamped;

    always @(*) begin
        if (current_money > 16'd10000)
            money_clamped = 16'd10000;
        else
            money_clamped = current_money;
    end

    //============================================================
    // 5�ڸ� ���� (��/õ/��/��/��)
    //============================================================
    reg [3:0] digit [0:4];  // digit[0] = ���� �ڸ�, digit[4] = ���� �ڸ�

    always @(*) begin
        digit[0] = (money_clamped / 10000) % 10;  // ��
        digit[1] = (money_clamped / 1000)  % 10;  // õ
        digit[2] = (money_clamped / 100)   % 10;  // ��
        digit[3] = (money_clamped / 10)    % 10;  // ��
        digit[4] = (money_clamped)         % 10;  // ��
    end

    //============================================================
    // �ڸ� ���� Multiplex Counter
    //============================================================
    reg [15:0] refresh_cnt = 0;
    reg [2:0]  digit_sel = 0;  // 0~4 �ݺ�

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            refresh_cnt <= 0;
            digit_sel   <= 0;
        end else begin
            refresh_cnt <= refresh_cnt + 1;

            // �� 1kHz ������ �ڸ� ���� (���� Ŭ�� 100MHz ����)
            if (refresh_cnt == 16'd2000) begin
                refresh_cnt <= 0;
                digit_sel <= (digit_sel == 4) ? 0 : digit_sel + 1;
            end
        end
    end

    //============================================================
    // ���� �� 7-seg ���� (active-low)
    //============================================================
    function [6:0] seg_decode;
        input [3:0] num;
        case(num)
            4'd0: seg_decode = ~7'b1000000;
            4'd1: seg_decode = ~7'b1111001;
            4'd2: seg_decode = ~7'b0100100;
            4'd3: seg_decode = ~7'b0110000;
            4'd4: seg_decode = ~7'b0011001;
            4'd5: seg_decode = ~7'b0010010;
            4'd6: seg_decode = ~7'b0000010;
            4'd7: seg_decode = ~7'b1111000;
            4'd8: seg_decode = ~7'b0000000;
            4'd9: seg_decode = ~7'b0010000;
            default: seg_decode = ~7'b1111111; // blank
        endcase
    endfunction

    //============================================================
    // Multiplex: digit_sel�� ���� an �� seg ����
    //============================================================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            an  <= 5'b11111;   // ��� ���� (active-low)
            seg <= 7'b1111111;
        end else begin
            case (digit_sel)
                0: begin  // ���� �ڸ�
                    an  <= 5'b01111;
                    seg <= seg_decode(digit[0]);
                end
                1: begin  // õ�� �ڸ�
                    an  <= 5'b10111;
                    seg <= seg_decode(digit[1]);
                end
                2: begin  // ���� �ڸ�
                    an  <= 5'b11011;
                    seg <= seg_decode(digit[2]);
                end
                3: begin  // ���� �ڸ�
                    an  <= 5'b11101;
                    seg <= seg_decode(digit[3]);
                end
                4: begin  // ���� �ڸ�
                    an  <= 5'b11110;
                    seg <= seg_decode(digit[4]);
                end
                default: begin
                    an  <= 5'b11111;
                    seg <= 7'b1111111;
                end
            endcase
        end
    end

endmodule
