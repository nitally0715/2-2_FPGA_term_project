//======================================================================
// Piezo_Buzzer.v (Rhythm FIXED Version)
// - ��ε� �ӵ��� ����� ���� �� �ִ� ���ڷ� ������
//======================================================================

module Piezo_Buzzer(
    input  wire clk,
    input  wire rst,

    input  wire [3:0] state,
    input  wire       spin_active,  // �귿�� ���� ȸ�� ���̸� 1
    input  wire       win_flag,     // �¸� ����

    output reg        piezo_out
);

    //==========================================================
    // FSM ���� ����
    //==========================================================
    localparam  S_IDLE         = 4'd0,
                S_BET_MONEY    = 4'd1,
                S_BET_SELECT   = 4'd2,
                S_NUMBER_INPUT = 4'd3,
                S_START_SPIN   = 4'd4,
                S_SLOW_DOWN    = 4'd5,
                S_STOP_RESULT  = 4'd6,
                S_WIN_DISPLAY  = 4'd7,
                S_LOSE_DISPLAY = 4'd8,
                S_UPDATE_MONEY = 4'd9,
                S_CHECK_MONEY  = 4'd10,
                S_NEXT_STAGE   = 4'd11,
                S_GAME_OVER    = 4'd12,
                S_GAME_CLEAR   = 4'd13;

    //==========================================================
    // �⺻ �� ���ļ� ����
    //==========================================================
    reg [31:0] tone_divider;
    reg [31:0] tone_cnt;
    reg        tone_clk;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            tone_cnt <= 0;
            tone_clk <= 0;
        end else begin
            if (tone_cnt >= tone_divider) begin
                tone_cnt <= 0;
                tone_clk <= ~tone_clk;
            end else begin
                tone_cnt <= tone_cnt + 1;
            end
        end
    end

    //==========================================================
    // ��ε� ����� ī����
    //==========================================================
    reg [31:0] mel_cnt;
    always @(posedge clk or posedge rst) begin
        if (rst)
            mel_cnt <= 0;
        else
            mel_cnt <= mel_cnt + 1;
    end

    //==========================================================
    // [����] ��Ʈ �ε����� ���� �����Ͽ� ���ڸ� ������ ����
    //==========================================================
    always @(*) begin
        case (state)

            //==================================================
            // �귿 ȸ���� (spin_active == 1)
            //==================================================
            S_START_SPIN, S_SLOW_DOWN: begin
                if (spin_active)
                    tone_divider = 32'd50000;   // 500Hz
                else
                    tone_divider = 32'd0;
            end

            //==================================================
            // �й��� : [25]�� ��Ʈ ��� (�� 0.67�� �ֱ� ������)
            //==================================================
            S_LOSE_DISPLAY: begin
                // [����] [20] -> [25] (�ӵ� ������)
                if ((mel_cnt[25] == 0)) 
                    tone_divider = 32'd90000;   // 277Hz (������)
                else
                    tone_divider = 32'd0;
            end

            //==================================================
            // �Ϲ� �¸� : [25:23] ��� (�� �ϳ��� �� 0.16��)
            // ��(0.16s) -> ��(0.16s) -> ��(0.16s) -> ����...
            //==================================================
            S_WIN_DISPLAY: begin
                // [����] [19:17] -> [25:23] (�ӵ� ������)
                case (mel_cnt[25:23])  
                    3'd0: tone_divider = 32'd35000;  // ��
                    3'd1: tone_divider = 32'd50000;  // ��
                    3'd2: tone_divider = 32'd70000;  // ��
                    default: tone_divider = 32'd0;   // ��� ����
                endcase
            end

            //==================================================
            // GAME_CLEAR : [26:24] ��� (�� �ϳ��� �� 0.33��)
            // õõ�� �����ϰ�
            //==================================================
            S_GAME_CLEAR: begin
                // [����] [21:19] -> [26:24] (�ӵ� ������)
                case (mel_cnt[26:24])
                    3'd0: tone_divider = 32'd30000; // A
                    3'd1: tone_divider = 32'd35000; // B
                    3'd2: tone_divider = 32'd30000; // A
                    3'd3: tone_divider = 32'd45000; // G
                    default: tone_divider = 32'd0;
                endcase
            end

            default: tone_divider = 0;
        endcase
    end

    //==========================================================
    // ���� piezo ��� (���� ó�� ����)
    //==========================================================
    always @(posedge clk or posedge rst) begin
        if (rst)
            piezo_out <= 0;
        else begin
            if (tone_divider == 0)
                piezo_out <= 0;
            else
                piezo_out <= tone_clk;
        end
    end

endmodule